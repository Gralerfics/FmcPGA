library IEEE;
use IEEE.std_logic_1164.all;

use work.types.all;


-- This module is used to accept resolved peripheral inputs and update the player state at a appropriate frequency.
entity player_state_updater is
    port (
        clk, rst: in std_logic
    );
end entity;


architecture Behavioral of player_state_updater is

begin

end architecture;
