library IEEE;
use IEEE.std_logic_1164.all;

use work.types.all;
use work.constants.all;


entity gamepad is
    -- port (
        
    -- );
end entity;


architecture Behavioral of gamepad is

begin

end architecture;
