library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.float_pkg.all;


entity top_module is

end entity;


architecture Behavioral of top_module is

begin

end architecture;
