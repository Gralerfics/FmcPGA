library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.numeric_std_unsigned.all;
use work.constants.all;


entity player_info is
    -- port (
        
    -- );
end entity;
