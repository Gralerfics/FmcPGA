library IEEE;
use IEEE.std_logic_1164.all;

use work.constants.all;


entity viewport_scanner is
    port (
        
    );
end entity;


architecture Behavioral of viewport_scanner is

begin

end architecture;
